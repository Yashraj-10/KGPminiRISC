`timescale 1ns/1ps

module alu_TB();
    //Inputs
    reg [31:0] a ;
    reg [31:0] b ;
    reg [3:0] ALUcntrl ;
    
    //Outputs
    wire [2:0] flag;
    wire [31:0] result;

    alu uut (
        .a(a),
        .b(b),
        .ALUcntrl(ALUcntrl),
        .flag(flag),
        .result(result)
    );

    initial begin 
        $monitor("time=%0d,a = %d, b = %d, ALUcntrl = %d, flag = %b, result = %d",$time, a, b, ALUcntrl, flag, result);
        #10 a = 32'b00000000000000000000000000000000; b = 32'b00000000000000000000000000000000; ALUcntrl = 4'b0000;
        #10 a = 32'b00000000000000000000000000000100; b = 32'b00000000000000000000000000000001; ALUcntrl = 4'b0000;
        #10 a = 32'b00000000000000000000000000000011; b = 32'b00000000000000000000000000000001; ALUcntrl = 4'b0001;
        #10 a = 32'b00000000000000000000000000000011; b = 32'b00000000000000000000000000000011; ALUcntrl = 4'b0010;
        #10 a = 32'b00000000000000000000000000000011; b = 32'b00000000000000000000000000000011; ALUcntrl = 4'b0011;
        #10 a = 32'b00000000000000000000000000000111; b = 32'b00000000000000000000000000000001; ALUcntrl = 4'b0101;
        #10 a = 32'b00000000000000000000000000000011; b = 32'b00000000000000000000000000000001; ALUcntrl = 4'b0110;
        #10 a = 32'b00000000000000000000000000001011; b = 32'b00000000000000000000000000000001; ALUcntrl = 4'b0111;
        #10 a = 32'b00000000000000000000000000001011; b = 32'b00000000000000000000000000100001; ALUcntrl = 4'b1000;
        #10 $finish;
    end
endmodule

